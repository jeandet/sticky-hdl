LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY bram_256x16 IS
    PORT (
        RDATA : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
        RADDR : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
        RCLK : IN STD_LOGIC;
        RCLKE : IN STD_LOGIC;
        RE : IN STD_LOGIC;
        WADDR : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
        WCLK : IN STD_LOGIC;
        WCLKE : IN STD_LOGIC;
        WDATA : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        MASK : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        WE : IN STD_LOGIC
    );
END ENTITY;

ARCHITECTURE hw_ram OF bram_256x16 IS
    COMPONENT SB_RAM40_4K
        GENERIC (
            INIT_0 : STRING;
            INIT_1 : STRING;
            INIT_2 : STRING;
            INIT_3 : STRING;
            INIT_4 : STRING;
            INIT_5 : STRING;
            INIT_6 : STRING;
            INIT_7 : STRING;
            INIT_8 : STRING;
            INIT_9 : STRING;
            INIT_A : STRING;
            INIT_B : STRING;
            INIT_C : STRING;
            INIT_D : STRING;
            INIT_E : STRING;
            INIT_F : STRING;
            READ_MODE : INTEGER;
            WRITE_MODE : INTEGER
        );
        PORT (
            RDATA : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
            RADDR : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
            RCLK : IN STD_LOGIC;
            RCLKE : IN STD_LOGIC;
            RE : IN STD_LOGIC;
            WADDR : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
            WCLK : IN STD_LOGIC;
            WCLKE : IN STD_LOGIC;
            WDATA : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
            MASK : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
            WE : IN STD_LOGIC
        );

    END COMPONENT;
BEGIN

    ram256x16_inst : SB_RAM40_4K GENERIC MAP(
        INIT_0 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_8 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_9 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_F => X"0000000000000000000000000000000000000000000000000000000000000000",
        READ_MODE => 0,
        WRITE_MODE => 0
    )
    PORT MAP(
        RDATA => RDATA,
        RADDR => "000" & RADDR,
        RCLK => RCLK,
        RCLKE => RCLKE,
        RE => RE,
        WADDR => "000" & WADDR,
        WCLK => WCLK,
        WCLKE => WCLKE,
        WDATA => WDATA,
        MASK => MASK,
        WE => WE
    );

END hw_ram;